module tb();

initial begin 
$display("a=%0d\n\tb=%0d\n\t\tc=%0d\n\t\t\td=%0d",10,20,30,40);
end

endmodule