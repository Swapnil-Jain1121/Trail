module tb();
#10;
endmodule
