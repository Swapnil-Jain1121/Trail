module tb();
#5;
endmodule
